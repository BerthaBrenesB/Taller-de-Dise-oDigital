library IEEE; use IEEE.STD_LOGIC_1164.all;
entity seven_seg_decoder is
	port(data: in STD_LOGIC_VECTOR(3 downto 0);
	segments: out STD_LOGIC_VECTOR(6 downto 0));
end;
architecture synth of seven_seg_decoder is
begin
	process(data) begin
		case data is
			--abcdefg
			when X"0" => segments <= "0000001";
			when X"1" => segments <= "1001111";
			when X"2" => segments <= "0010010";
			when X"3" => segments <= "0000110";
			when X"4" => segments <= "1001100";
			when X"5" => segments <= "0100100";
			when X"6" => segments <= "0100000";
			when X"7" => segments <= "0001111";
			when X"8" => segments <= "0000000";
			when X"9" => segments <= "0000100";
			when others => segments <= "0000000";
		end case;
	end process;
end;